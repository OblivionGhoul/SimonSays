module Tone_Generator (
    input  logic        clk,
    input  logic        rst,
    input  logic [9:0]  frequency,       // Frequency in Hz (0 = silence)
    input  logic [15:0] ticks_per_milli, // Ticks per millisecond for timing
    output logic        sound            // Output tone signal
);

    logic [31:0] tick_counter;
    logic [31:0] ticks_per_second;

    assign ticks_per_second = ticks_per_milli * 1000; // Calculate ticks per second

    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            tick_counter <= 0;
            sound <= 0;
        end else if (frequency == 0) begin
            sound <= 0; // Silence when frequency is 0
        end else begin
            tick_counter <= tick_counter + frequency; // Increment by the frequency
            if (tick_counter >= (ticks_per_second >> 1)) begin
                sound <= ~sound; // Toggle sound signal
                tick_counter <= tick_counter - (ticks_per_second >> 1);
            end
        end
    end

endmodule
